module complement (
    input clk,
    input rst,
    input clr,
    input data_in,
    output reg data_out
);

reg d;

always@(posedge clk) begin
    if (rst || clr) begin
        data_out <= 1'b0;
        d <= 1'b0;
    end else begin
        data_out <= d ^ data_in; // XOR operation
        d <= d | data_in; // OR operation
    end
end
    
endmodule